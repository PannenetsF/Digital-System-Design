$date
	Tue Dec  1 09:14:10 2020
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module test $end
$var wire 10 ! LEDR [9:0] $end
$var reg 1 " CLOCK_50 $end
$var reg 1 # KEY $end
$var reg 2 $ SW [1:0] $end
$scope module u $end
$var wire 1 " CLOCK_50 $end
$var wire 1 # KEY [2:2] $end
$var wire 10 % LEDR [9:0] $end
$var wire 2 & SW [17:16] $end
$var wire 1 ' reset $end
$var wire 1 ( push $end
$var wire 1 ) en $end
$var wire 1 * clk $end
$var reg 2 + cnt [1:0] $end
$var reg 10 , f_0_to_9 [9:0] $end
$var reg 10 - f_9_to_0 [9:0] $end
$var reg 1 . read $end
$var reg 4 / timer [3:0] $end
$scope module u_sync $end
$var wire 1 . read $end
$var wire 1 ' reset $end
$var wire 1 # sig $end
$var wire 1 * clk $end
$var reg 1 0 sig_buf $end
$var reg 1 ( valid $end
$upscope $end
$scope module u_tik $end
$var wire 1 " CLOCK_50 $end
$var wire 1 ' reset $end
$var reg 32 1 cnt [31:0] $end
$var reg 1 * tik $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
bx 1
00
bx /
x.
bx -
bx ,
bx +
x*
x)
x(
x'
bx &
bx %
bx $
0#
0"
bx !
$end
#1
b0 !
b0 %
0(
b0 /
0.
b0 +
b0 -
b0 ,
0*
b0 1
1'
b1x $
b1x &
1"
#2
1)
0'
b1 $
b1 &
0"
#3
b1 1
1"
#4
0"
#5
b10 1
1"
#6
0"
#7
b11 1
1"
#8
0"
#9
b100 1
1"
#10
0"
#11
b101 1
1"
#12
0"
#13
b110 1
1"
#14
0"
#15
b111 1
1"
#16
0"
#17
b1000 1
1"
#18
0"
#19
b1001 1
1"
#20
0"
#21
b1010 1
1"
#22
0"
#23
b1011 1
1"
#24
0"
#25
b1100 1
1"
#26
0"
#27
b1101 1
1"
#28
0"
#29
b1110 1
1"
#30
0"
#31
b1111 1
1"
#32
0"
#33
b10000 1
1"
#34
0"
#35
b10001 1
1"
#36
0"
#37
b10010 1
1"
#38
0"
#39
b10011 1
1"
#40
0"
#41
b10100 1
1"
#42
0"
#43
b10101 1
1"
#44
0"
#45
b10110 1
1"
#46
0"
#47
b10111 1
1"
#48
0"
#49
b11000 1
1"
#50
0"
#51
b11001 1
1"
#52
0"
#53
b11010 1
1"
#54
0"
#55
b11011 1
1"
#56
0"
#57
b11100 1
1"
#58
0"
#59
b11101 1
1"
#60
0"
#61
b11110 1
1"
#62
10
0"
1#
#63
b11111 1
00
1"
0#
#64
0"
#65
b100000 1
1"
#66
0"
#67
b100001 1
1"
#68
0"
#69
b100010 1
1"
#70
0"
#71
b100011 1
1"
#72
0"
#73
b100100 1
1"
#74
0"
#75
b100101 1
1"
#76
0"
#77
b100110 1
1"
#78
0"
#79
b100111 1
1"
#80
0"
#81
b101000 1
1"
#82
0"
#83
b101001 1
1"
#84
0"
#85
b101010 1
1"
#86
0"
#87
b101011 1
1"
#88
0"
#89
b101100 1
1"
#90
0"
#91
b101101 1
1"
#92
0"
#93
b101110 1
1"
#94
0"
#95
b101111 1
1"
#96
0"
#97
b110000 1
1"
#98
0"
#99
b110001 1
1"
#100
0"
#101
b110010 1
1"
#102
0"
#103
b110011 1
1"
#104
0"
#105
b110100 1
1"
#106
0"
#107
b110101 1
1"
#108
0"
#109
b110110 1
1"
#110
0"
#111
b110111 1
1"
#112
0"
#113
b111000 1
1"
#114
0"
#115
b111001 1
1"
#116
0"
#117
b111010 1
1"
#118
0"
#119
b111011 1
1"
#120
0"
#121
b111100 1
1"
#122
0"
#123
b111101 1
10
1"
1#
#124
00
0"
0#
#125
b111110 1
1"
#126
0"
#127
b111111 1
1"
#128
0"
#129
b1000000 1
1"
#130
0"
#131
b1000001 1
1"
#132
0"
#133
b1000010 1
1"
#134
0"
#135
b1000011 1
1"
#136
0"
#137
b1000100 1
1"
#138
0"
#139
b1000101 1
1"
#140
0"
#141
b1000110 1
1"
#142
0"
#143
b1000111 1
1"
#144
0"
#145
b1001000 1
1"
#146
0"
#147
b1001001 1
1"
#148
0"
#149
b1001010 1
1"
#150
0"
#151
b1001011 1
1"
#152
0"
#153
b1001100 1
1"
#154
0"
#155
b1001101 1
1"
#156
0"
#157
b1001110 1
1"
#158
0"
#159
b1001111 1
1"
#160
0"
#161
b1010000 1
1"
#162
0"
#163
b1010001 1
1"
#164
0"
#165
b1010010 1
1"
#166
0"
#167
b1010011 1
1"
#168
0"
#169
b1010100 1
1"
#170
0"
#171
b1010101 1
1"
#172
0"
#173
b1010110 1
1"
#174
0"
#175
b1010111 1
1"
#176
0"
#177
b1011000 1
1"
#178
0"
#179
b1011001 1
1"
#180
0"
#181
b1011010 1
1"
#182
0"
#183
b1011011 1
1"
#184
10
0"
1#
#185
b1011100 1
00
1"
0#
#186
0"
#187
b1011101 1
1"
#188
0"
#189
b1011110 1
1"
#190
0"
#191
b1011111 1
1"
#192
0"
#193
b1100000 1
1"
#194
0"
#195
b1100001 1
1"
#196
0"
#197
b1100010 1
1"
#198
0"
#199
b1100011 1
1"
#200
0"
#201
b1100100 1
1"
#202
0"
#203
b1100101 1
1"
#204
0"
#205
b1100110 1
1"
#206
0"
#207
b1100111 1
1"
#208
0"
#209
b1101000 1
1"
#210
0"
#211
b1101001 1
1"
#212
0"
#213
b1101010 1
1"
#214
0"
#215
b1101011 1
1"
#216
0"
#217
b1101100 1
1"
#218
0"
#219
b1101101 1
1"
#220
0"
#221
b1101110 1
1"
#222
0"
#223
b1101111 1
1"
#224
0"
#225
b1110000 1
1"
#226
0"
#227
b1110001 1
1"
#228
0"
#229
b1110010 1
1"
#230
0"
#231
b1110011 1
1"
#232
0"
#233
b1110100 1
1"
#234
0"
#235
b1110101 1
1"
#236
0"
#237
b1110110 1
1"
#238
0"
#239
b1110111 1
1"
#240
0"
#241
b1111000 1
1"
#242
0"
#243
b1111001 1
1"
#244
0"
#245
b1111010 1
1"
#246
0"
#247
b1111011 1
1"
#248
0"
#249
b1111100 1
1"
#250
0"
#251
b1111101 1
1"
#252
0"
#253
b1111110 1
1"
#254
0"
#255
b1111111 1
1"
#256
0"
#257
b10000000 1
1"
#258
0"
#259
b10000001 1
1"
#260
0"
#261
b10000010 1
1"
#262
0"
#263
b10000011 1
1"
#264
0"
#265
b10000100 1
1"
#266
0"
#267
b10000101 1
1"
#268
0"
#269
b10000110 1
1"
#270
0"
#271
b10000111 1
1"
#272
0"
#273
b10001000 1
1"
#274
0"
#275
b10001001 1
1"
#276
0"
#277
b10001010 1
1"
#278
0"
#279
b10001011 1
1"
#280
0"
#281
b10001100 1
1"
#282
0"
#283
b10001101 1
1"
#284
0"
#285
b10001110 1
1"
#286
0"
#287
b10001111 1
1"
#288
0"
#289
b10010000 1
1"
#290
0"
#291
b10010001 1
1"
#292
0"
#293
b10010010 1
1"
#294
0"
#295
b10010011 1
1"
#296
0"
#297
b10010100 1
1"
#298
0"
#299
b10010101 1
1"
#300
0"
#301
b10010110 1
1"
#302
0"
#303
b10010111 1
1"
#304
0"
#305
b10011000 1
1"
#306
0"
#307
b10011001 1
1"
#308
0"
#309
b10011010 1
1"
#310
0"
#311
b10011011 1
1"
#312
0"
#313
b10011100 1
1"
#314
0"
#315
b10011101 1
1"
#316
0"
#317
b10011110 1
1"
#318
0"
#319
b10011111 1
1"
#320
0"
#321
b10100000 1
1"
#322
0"
#323
b10100001 1
1"
#324
0"
#325
b10100010 1
1"
#326
0"
#327
b10100011 1
1"
#328
0"
#329
b10100100 1
1"
#330
0"
#331
b10100101 1
1"
#332
0"
#333
b10100110 1
1"
#334
0"
#335
b10100111 1
1"
#336
0"
#337
b10101000 1
1"
#338
0"
#339
b10101001 1
1"
#340
0"
#341
b10101010 1
1"
#342
0"
#343
b10101011 1
1"
#344
0"
#345
b10101100 1
1"
#346
0"
#347
b10101101 1
1"
#348
0"
#349
b10101110 1
1"
#350
0"
#351
b10101111 1
1"
#352
0"
#353
b10110000 1
1"
#354
0"
#355
b10110001 1
1"
#356
0"
#357
b10110010 1
1"
#358
0"
#359
b10110011 1
1"
#360
0"
#361
b10110100 1
1"
#362
0"
#363
b10110101 1
1"
#364
0"
#365
b10110110 1
1"
#366
0"
#367
b10110111 1
1"
#368
0"
#369
b10111000 1
1"
#370
0"
#371
b10111001 1
1"
#372
0"
#373
b10111010 1
1"
#374
0"
#375
b10111011 1
1"
#376
0"
#377
b10111100 1
1"
#378
0"
#379
b10111101 1
1"
#380
0"
#381
b10111110 1
1"
#382
0"
#383
b10111111 1
1"
#384
0"
#385
b11000000 1
1"
